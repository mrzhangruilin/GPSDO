module Preheat(
    input   CLK_Sys,            //系统10M时钟
    input   CLK_Rst,            //复位信号

    output  Flag_Preheat_Done    //预热完成标志位
);





endmodule
